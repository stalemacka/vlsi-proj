entity cpu is
end cpu;