entity cpu is
