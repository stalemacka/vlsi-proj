library ieee;
use ieee.std_logic_1164.all;

entity cpu is
port(abus: std_logic_vector(31 downto 0));
end cpu;

architecture cpu_behav of cpu is
begin
end cpu_behav;